`timescale 1ns/1ns
module tb_LED_7_Thanh;
//testbench body
parameter N= ;
parameter END_TIME=100;
parameter VALUE_NUM=2*N;



endmodule